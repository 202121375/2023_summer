module fifo(
    clk,
    n_rst,
    tx_data,
    rx_data,
    rx_fifo,
    result
);

    input clk;
    input n_rst;
    output tx_data;
    output rx_fifo;

    
endmodule